// n=32 w=16               


module APPR (AH,AL,BH,BL,PP1,carry);
	input [15:0]AH,BH,AL,BL;
	output [14:0]PP1;
	output carry;
	wire P0,P1,P2,P3,P4,P5,P6,P7,O0,O1,O2,O3,O4,O5,O6,O7;

	assign P0=(BL[1]&AH[15])|(BL[2]&AH[14])|(BL[3]&AH[13])|(BL[4]&AH[12])|(BL[5]&AH[11])|(BL[6]&AH[10])|(BL[7]&AH[9])|(BL[8]&AH[8])|(BL[9]&AH[7])|(BL[10]&AH[6])|(BL[11]&AH[5])|(BL[12]&AH[4])|(BL[13]&AH[3])|(BL[14]&AH[2])|(BL[15]&AH[1]);
	assign P1=(BL[2]&AH[15])|(BL[3]&AH[14])|(BL[4]&AH[13])|(BL[5]&AH[12])|(BL[6]&AH[11])|(BL[7]&AH[10])|(BL[8]&AH[9])|(BL[9]&AH[8])|(BL[10]&AH[7])|(BL[11]&AH[6])|(BL[12]&AH[5])|(BL[13]&AH[4])|(BL[14]&AH[3])|(BL[15]&AH[2]);
	assign P2=(BL[3]&AH[15])|(BL[4]&AH[14])|(BL[5]&AH[13])|(BL[6]&AH[12])|(BL[7]&AH[11])|(BL[8]&AH[10])|(BL[9]&AH[9])|(BL[10]&AH[8])|(BL[11]&AH[7])|(BL[12]&AH[6])|(BL[13]&AH[5])|(BL[14]&AH[4])|(BL[15]&AH[3]);
	assign P3=(BL[4]&AH[15])|(BL[5]&AH[14])|(BL[6]&AH[13])|(BL[7]&AH[12])|(BL[8]&AH[11])|(BL[9]&AH[10])|(BL[10]&AH[9])|(BL[11]&AH[8])|(BL[12]&AH[7])|(BL[13]&AH[6])|(BL[14]&AH[5])|(BL[15]&AH[4]);
	assign P4=(BL[5]&AH[15])|(BL[6]&AH[14])|(BL[7]&AH[13])|(BL[8]&AH[12])|(BL[9]&AH[11])|(BL[10]&AH[10])|(BL[11]&AH[9])|(BL[12]&AH[8])|(BL[13]&AH[7])|(BL[14]&AH[6])|(BL[15]&AH[5]);
	assign P5=(BL[6]&AH[15])|(BL[7]&AH[14])|(BL[8]&AH[13])|(BL[9]&AH[12])|(BL[10]&AH[11])|(BL[11]&AH[10])|(BL[12]&AH[9])|(BL[13]&AH[8])|(BL[14]&AH[7])|(BL[15]&AH[6]);
	assign P6=(BL[7]&AH[15])|(BL[8]&AH[14])|(BL[9]&AH[13])|(BL[10]&AH[12])|(BL[11]&AH[11])|(BL[12]&AH[10])|(BL[13]&AH[9])|(BL[14]&AH[8])|(BL[15]&AH[7]);
	assign P7=(BL[8]&AH[15])|(BL[9]&AH[14])|(BL[10]&AH[13])|(BL[11]&AH[12])|(BL[12]&AH[11])|(BL[13]&AH[10])|(BL[14]&AH[9])|(BL[15]&AH[8]);
	assign P8=(BL[9]&AH[15])|(BL[10]&AH[14])|(BL[11]&AH[13])|(BL[12]&AH[12])|(BL[13]&AH[11])|(BL[14]&AH[10])|(BL[15]&AH[9]);
	assign P9=(BL[10]&AH[15])|(BL[11]&AH[14])|(BL[12]&AH[13])|(BL[13]&AH[12])|(BL[14]&AH[11])|(BL[15]&AH[10]);
	assign P10=(BL[11]&AH[15])|(BL[12]&AH[14])|(BL[13]&AH[13])|(BL[14]&AH[12])|(BL[15]&AH[11]);
	assign P11=(BL[12]&AH[15])|(BL[13]&AH[14])|(BL[14]&AH[13])|(BL[15]&AH[12]);
	assign P12=(BL[13]&AH[15])|(BL[14]&AH[14])|(BL[15]&AH[13]);
	assign P13=(BL[14]&AH[15])|(BL[15]&AH[14]);
	assign P14=(BL[15]&AH[15]);
	assign P15=P14&P13;
	assign O0=(AL[1]&BH[15])|(AL[2]&BH[14])|(AL[3]&BH[13])|(AL[4]&BH[12])|(AL[5]&BH[11])|(AL[6]&BH[10])|(AL[7]&BH[9])|(AL[8]&BH[8])|(AL[9]&BH[7])|(AL[10]&BH[6])|(AL[11]&BH[5])|(AL[12]&BH[4])|(AL[13]&BH[3])|(AL[14]&BH[2])|(AL[15]&BH[1]);
	assign O1=(AL[2]&BH[15])|(AL[3]&BH[14])|(AL[4]&BH[13])|(AL[5]&BH[12])|(AL[6]&BH[11])|(AL[7]&BH[10])|(AL[8]&BH[9])|(AL[9]&BH[8])|(AL[10]&BH[7])|(AL[11]&BH[6])|(AL[12]&BH[5])|(AL[13]&BH[4])|(AL[14]&BH[3])|(AL[15]&BH[2]);
	assign O2=(AL[3]&BH[15])|(AL[4]&BH[14])|(AL[5]&BH[13])|(AL[6]&BH[12])|(AL[7]&BH[11])|(AL[8]&BH[10])|(AL[9]&BH[9])|(AL[10]&BH[8])|(AL[11]&BH[7])|(AL[12]&BH[6])|(AL[13]&BH[5])|(AL[14]&BH[4])|(AL[15]&BH[3]);
	assign O3=(AL[4]&BH[15])|(AL[5]&BH[14])|(AL[6]&BH[13])|(AL[7]&BH[12])|(AL[8]&BH[11])|(AL[9]&BH[10])|(AL[10]&BH[9])|(AL[11]&BH[8])|(AL[12]&BH[7])|(AL[13]&BH[6])|(AL[14]&BH[5])|(AL[15]&BH[4]);
	assign O4=(AL[5]&BH[15])|(AL[6]&BH[14])|(AL[7]&BH[13])|(AL[8]&BH[12])|(AL[9]&BH[11])|(AL[10]&BH[10])|(AL[11]&BH[9])|(AL[12]&BH[8])|(AL[13]&BH[7])|(AL[14]&BH[6])|(AL[15]&BH[5]);
	assign O5=(AL[6]&BH[15])|(AL[7]&BH[14])|(AL[8]&BH[13])|(AL[9]&BH[12])|(AL[10]&BH[11])|(AL[11]&BH[10])|(AL[12]&BH[9])|(AL[13]&BH[8])|(AL[14]&BH[7])|(AL[15]&BH[6]);
	assign O6=(AL[7]&BH[15])|(AL[8]&BH[14])|(AL[9]&BH[13])|(AL[10]&BH[12])|(AL[11]&BH[11])|(AL[12]&BH[10])|(AL[13]&BH[9])|(AL[14]&BH[8])|(AL[15]&BH[7]);
	assign O7=(AL[8]&BH[15])|(AL[9]&BH[14])|(AL[10]&BH[13])|(AL[11]&BH[12])|(AL[12]&BH[11])|(AL[13]&BH[10])|(AL[14]&BH[9])|(AL[15]&BH[8]);
	assign O8=(AL[9]&BH[15])|(AL[10]&BH[14])|(AL[11]&BH[13])|(AL[12]&BH[12])|(AL[13]&BH[11])|(AL[14]&BH[10])|(AL[15]&BH[9]);
	assign O9=(AL[10]&BH[15])|(AL[11]&BH[14])|(AL[12]&BH[13])|(AL[13]&BH[12])|(AL[14]&BH[11])|(AL[15]&BH[10]);
	assign O10=(AL[11]&BH[15])|(AL[12]&BH[14])|(AL[13]&BH[13])|(AL[14]&BH[12])|(AL[15]&BH[11]);
	assign O11=(AL[12]&BH[15])|(AL[13]&BH[14])|(AL[14]&BH[13])|(AL[15]&BH[12]);
	assign O12=(AL[13]&BH[15])|(AL[14]&BH[14])|(AL[15]&BH[13]);
	assign O13=(AL[14]&BH[15])|(AL[15]&BH[14]);
	assign O14=(AL[15]&BH[15]);
	assign O15=O14&O13;
	assign PP1[0]=P0|O0;
	assign PP1[1]=P1|O1;
	assign PP1[2]=P2|O2;
	assign PP1[3]=P3|O3;
	assign PP1[4]=P4|O4;
	assign PP1[5]=P5|O5;
	assign PP1[6]=P6|O6;
	assign PP1[7]=P7|O7;
	assign PP1[8]=P8|O8;
	assign PP1[9]=P9|O9;
	assign PP1[10]=P10|O10;
	assign PP1[11]=P11|O11;
	assign PP1[12]=P12|O12;
	assign PP1[13]=P13|O13;
	assign PP1[14]=P14|O14;
	assign carry= P15|O15;
endmodule

//******************* LSD ***************************
module LSD_n32_ss16(X,Kx,XH,XL);
	input [31:0]X;
	output Kx;
	output [15:0]XH;
	output [15:0]XL;
	assign Kx=(X[31] | X[30] | X[29] | X[28] | X[27] | X[26] | X[25] | X[24]|X[23] | X[22] | X[21] | X[20] | X[19] | X[18] | X[17] | X[16]) ? 1'b1:1'b0;

	assign XH=(Kx==1'b1) ? X[31:16]:X[15:0];

	assign XL=(Kx==1'b1) ? X[15:0]:16'b0;
endmodule
//**********************HA and FA***********************
module HA(A,B,sum,carry);
    input A, B;
    output sum, carry;
	assign sum = A ^ B;   // XOR operation for sum
	assign carry = A & B; // AND operation for carry
endmodule


module FA (A,B,cin,sum,cout);
    input A, B, cin;
    output sum, cout;
	assign sum = A ^ B ^ cin;
	assign cout = (A & B) | (cin & (A ^ B));
endmodule






//******************* wallace 4 ***************************
module wallace_with_carry(A,B,carry,FinalOut_MSB,FinalOut_LSB);
input [15:0]A,B;
input carry;
output [16:0]FinalOut_MSB;
output [14:0]FinalOut_LSB;
wire [31:0] FinalOut;

//**************************************Generating PPs**************
assign FinalOut[0]=A[0] & B[0];
assign OL0X1C1= A[1] & B[0];
assign OL0X2C1= A[0] & B[1];
assign OL0X1C2= A[2] & B[0];
assign OL0X2C2= A[1] & B[1];
assign OL0X3C2= A[0] & B[2];
assign OL0X1C3= A[3] & B[0];
assign OL0X2C3= A[2] & B[1];
assign OL0X3C3= A[1] & B[2];
assign OL0X4C3= A[0] & B[3];
assign OL0X1C4= A[4] & B[0];
assign OL0X2C4= A[3] & B[1];
assign OL0X3C4= A[2] & B[2];
assign OL0X4C4= A[1] & B[3];
assign OL0X5C4= A[0] & B[4];
assign OL0X1C5= A[5] & B[0];
assign OL0X2C5= A[4] & B[1];
assign OL0X3C5= A[3] & B[2];
assign OL0X4C5= A[2] & B[3];
assign OL0X5C5= A[1] & B[4];
assign OL0X6C5= A[0] & B[5];
assign OL0X1C6= A[6] & B[0];
assign OL0X2C6= A[5] & B[1];
assign OL0X3C6= A[4] & B[2];
assign OL0X4C6= A[3] & B[3];
assign OL0X5C6= A[2] & B[4];
assign OL0X6C6= A[1] & B[5];
assign OL0X7C6= A[0] & B[6];
assign OL0X1C7= A[7] & B[0];
assign OL0X2C7= A[6] & B[1];
assign OL0X3C7= A[5] & B[2];
assign OL0X4C7= A[4] & B[3];
assign OL0X5C7= A[3] & B[4];
assign OL0X6C7= A[2] & B[5];
assign OL0X7C7= A[1] & B[6];
assign OL0X8C7= A[0] & B[7];
assign OL0X1C8= A[8] & B[0];
assign OL0X2C8= A[7] & B[1];
assign OL0X3C8= A[6] & B[2];
assign OL0X4C8= A[5] & B[3];
assign OL0X5C8= A[4] & B[4];
assign OL0X6C8= A[3] & B[5];
assign OL0X7C8= A[2] & B[6];
assign OL0X8C8= A[1] & B[7];
assign OL0X9C8= A[0] & B[8];
assign OL0X1C9= A[9] & B[0];
assign OL0X2C9= A[8] & B[1];
assign OL0X3C9= A[7] & B[2];
assign OL0X4C9= A[6] & B[3];
assign OL0X5C9= A[5] & B[4];
assign OL0X6C9= A[4] & B[5];
assign OL0X7C9= A[3] & B[6];
assign OL0X8C9= A[2] & B[7];
assign OL0X9C9= A[1] & B[8];
assign OL0X10C9= A[0] & B[9];
assign OL0X1C10= A[10] & B[0];
assign OL0X2C10= A[9] & B[1];
assign OL0X3C10= A[8] & B[2];
assign OL0X4C10= A[7] & B[3];
assign OL0X5C10= A[6] & B[4];
assign OL0X6C10= A[5] & B[5];
assign OL0X7C10= A[4] & B[6];
assign OL0X8C10= A[3] & B[7];
assign OL0X9C10= A[2] & B[8];
assign OL0X10C10= A[1] & B[9];
assign OL0X11C10= A[0] & B[10];
assign OL0X1C11= A[11] & B[0];
assign OL0X2C11= A[10] & B[1];
assign OL0X3C11= A[9] & B[2];
assign OL0X4C11= A[8] & B[3];
assign OL0X5C11= A[7] & B[4];
assign OL0X6C11= A[6] & B[5];
assign OL0X7C11= A[5] & B[6];
assign OL0X8C11= A[4] & B[7];
assign OL0X9C11= A[3] & B[8];
assign OL0X10C11= A[2] & B[9];
assign OL0X11C11= A[1] & B[10];
assign OL0X12C11= A[0] & B[11];
assign OL0X1C12= A[12] & B[0];
assign OL0X2C12= A[11] & B[1];
assign OL0X3C12= A[10] & B[2];
assign OL0X4C12= A[9] & B[3];
assign OL0X5C12= A[8] & B[4];
assign OL0X6C12= A[7] & B[5];
assign OL0X7C12= A[6] & B[6];
assign OL0X8C12= A[5] & B[7];
assign OL0X9C12= A[4] & B[8];
assign OL0X10C12= A[3] & B[9];
assign OL0X11C12= A[2] & B[10];
assign OL0X12C12= A[1] & B[11];
assign OL0X13C12= A[0] & B[12];
assign OL0X1C13= A[13] & B[0];
assign OL0X2C13= A[12] & B[1];
assign OL0X3C13= A[11] & B[2];
assign OL0X4C13= A[10] & B[3];
assign OL0X5C13= A[9] & B[4];
assign OL0X6C13= A[8] & B[5];
assign OL0X7C13= A[7] & B[6];
assign OL0X8C13= A[6] & B[7];
assign OL0X9C13= A[5] & B[8];
assign OL0X10C13= A[4] & B[9];
assign OL0X11C13= A[3] & B[10];
assign OL0X12C13= A[2] & B[11];
assign OL0X13C13= A[1] & B[12];
assign OL0X14C13= A[0] & B[13];
assign OL0X1C14= A[14] & B[0];
assign OL0X2C14= A[13] & B[1];
assign OL0X3C14= A[12] & B[2];
assign OL0X4C14= A[11] & B[3];
assign OL0X5C14= A[10] & B[4];
assign OL0X6C14= A[9] & B[5];
assign OL0X7C14= A[8] & B[6];
assign OL0X8C14= A[7] & B[7];
assign OL0X9C14= A[6] & B[8];
assign OL0X10C14= A[5] & B[9];
assign OL0X11C14= A[4] & B[10];
assign OL0X12C14= A[3] & B[11];
assign OL0X13C14= A[2] & B[12];
assign OL0X14C14= A[1] & B[13];
assign OL0X15C14= A[0] & B[14];
//************************for (n-1)th Column*************
assign OL0X1C15= A[15] & B[0];
assign OL0X2C15= A[14] & B[1];
assign OL0X3C15= A[13] & B[2];
assign OL0X4C15= A[12] & B[3];
assign OL0X5C15= A[11] & B[4];
assign OL0X6C15= A[10] & B[5];
assign OL0X7C15= A[9] & B[6];
assign OL0X8C15= A[8] & B[7];
assign OL0X9C15= A[7] & B[8];
assign OL0X10C15= A[6] & B[9];
assign OL0X11C15= A[5] & B[10];
assign OL0X12C15= A[4] & B[11];
assign OL0X13C15= A[3] & B[12];
assign OL0X14C15= A[2] & B[13];
assign OL0X15C15= A[1] & B[14];
assign OL0X16C15= A[0] & B[15];
//************************for (n)th Column*************
assign OL0X1C16= A[15] & B[1];
assign OL0X2C16= A[14] & B[2];
assign OL0X3C16= A[13] & B[3];
assign OL0X4C16= A[12] & B[4];
assign OL0X5C16= A[11] & B[5];
assign OL0X6C16= A[10] & B[6];
assign OL0X7C16= A[9] & B[7];
assign OL0X8C16= A[8] & B[8];
assign OL0X9C16= A[7] & B[9];
assign OL0X10C16= A[6] & B[10];
assign OL0X11C16= A[5] & B[11];
assign OL0X12C16= A[4] & B[12];
assign OL0X13C16= A[3] & B[13];
assign OL0X14C16= A[2] & B[14];
assign OL0X15C16= A[1] & B[15];
//******************************for the rest of Columns except for the last one************
assign OL0X1C17= A[15] & B[2];
assign OL0X2C17= A[14] & B[3];
assign OL0X3C17= A[13] & B[4];
assign OL0X4C17= A[12] & B[5];
assign OL0X5C17= A[11] & B[6];
assign OL0X6C17= A[10] & B[7];
assign OL0X7C17= A[9] & B[8];
assign OL0X8C17= A[8] & B[9];
assign OL0X9C17= A[7] & B[10];
assign OL0X10C17= A[6] & B[11];
assign OL0X11C17= A[5] & B[12];
assign OL0X12C17= A[4] & B[13];
assign OL0X13C17= A[3] & B[14];
assign OL0X14C17= A[2] & B[15];
assign OL0X1C18= A[15] & B[3];
assign OL0X2C18= A[14] & B[4];
assign OL0X3C18= A[13] & B[5];
assign OL0X4C18= A[12] & B[6];
assign OL0X5C18= A[11] & B[7];
assign OL0X6C18= A[10] & B[8];
assign OL0X7C18= A[9] & B[9];
assign OL0X8C18= A[8] & B[10];
assign OL0X9C18= A[7] & B[11];
assign OL0X10C18= A[6] & B[12];
assign OL0X11C18= A[5] & B[13];
assign OL0X12C18= A[4] & B[14];
assign OL0X13C18= A[3] & B[15];
assign OL0X1C19= A[15] & B[4];
assign OL0X2C19= A[14] & B[5];
assign OL0X3C19= A[13] & B[6];
assign OL0X4C19= A[12] & B[7];
assign OL0X5C19= A[11] & B[8];
assign OL0X6C19= A[10] & B[9];
assign OL0X7C19= A[9] & B[10];
assign OL0X8C19= A[8] & B[11];
assign OL0X9C19= A[7] & B[12];
assign OL0X10C19= A[6] & B[13];
assign OL0X11C19= A[5] & B[14];
assign OL0X12C19= A[4] & B[15];
assign OL0X1C20= A[15] & B[5];
assign OL0X2C20= A[14] & B[6];
assign OL0X3C20= A[13] & B[7];
assign OL0X4C20= A[12] & B[8];
assign OL0X5C20= A[11] & B[9];
assign OL0X6C20= A[10] & B[10];
assign OL0X7C20= A[9] & B[11];
assign OL0X8C20= A[8] & B[12];
assign OL0X9C20= A[7] & B[13];
assign OL0X10C20= A[6] & B[14];
assign OL0X11C20= A[5] & B[15];
assign OL0X1C21= A[15] & B[6];
assign OL0X2C21= A[14] & B[7];
assign OL0X3C21= A[13] & B[8];
assign OL0X4C21= A[12] & B[9];
assign OL0X5C21= A[11] & B[10];
assign OL0X6C21= A[10] & B[11];
assign OL0X7C21= A[9] & B[12];
assign OL0X8C21= A[8] & B[13];
assign OL0X9C21= A[7] & B[14];
assign OL0X10C21= A[6] & B[15];
assign OL0X1C22= A[15] & B[7];
assign OL0X2C22= A[14] & B[8];
assign OL0X3C22= A[13] & B[9];
assign OL0X4C22= A[12] & B[10];
assign OL0X5C22= A[11] & B[11];
assign OL0X6C22= A[10] & B[12];
assign OL0X7C22= A[9] & B[13];
assign OL0X8C22= A[8] & B[14];
assign OL0X9C22= A[7] & B[15];
assign OL0X1C23= A[15] & B[8];
assign OL0X2C23= A[14] & B[9];
assign OL0X3C23= A[13] & B[10];
assign OL0X4C23= A[12] & B[11];
assign OL0X5C23= A[11] & B[12];
assign OL0X6C23= A[10] & B[13];
assign OL0X7C23= A[9] & B[14];
assign OL0X8C23= A[8] & B[15];
assign OL0X1C24= A[15] & B[9];
assign OL0X2C24= A[14] & B[10];
assign OL0X3C24= A[13] & B[11];
assign OL0X4C24= A[12] & B[12];
assign OL0X5C24= A[11] & B[13];
assign OL0X6C24= A[10] & B[14];
assign OL0X7C24= A[9] & B[15];
assign OL0X1C25= A[15] & B[10];
assign OL0X2C25= A[14] & B[11];
assign OL0X3C25= A[13] & B[12];
assign OL0X4C25= A[12] & B[13];
assign OL0X5C25= A[11] & B[14];
assign OL0X6C25= A[10] & B[15];
assign OL0X1C26= A[15] & B[11];
assign OL0X2C26= A[14] & B[12];
assign OL0X3C26= A[13] & B[13];
assign OL0X4C26= A[12] & B[14];
assign OL0X5C26= A[11] & B[15];
assign OL0X1C27= A[15] & B[12];
assign OL0X2C27= A[14] & B[13];
assign OL0X3C27= A[13] & B[14];
assign OL0X4C27= A[12] & B[15];
assign OL0X1C28= A[15] & B[13];
assign OL0X2C28= A[14] & B[14];
assign OL0X3C28= A[13] & B[15];
assign OL0X1C29= A[15] & B[14];
assign OL0X2C29= A[14] & B[15];
//*******************************for the last column of PPS*****************
assign OL0X1C30= A[15] & B[15];
//*********************************************END of Generating Partial Products********************************************************
//***********************************Begin of Level 1 ************************************
assign {OL1X1C2,FinalOut[1]}=OL0X2C1+OL0X1C1;
assign {OL1X1C3,OL1X2C2}=OL0X3C2+OL0X2C2+OL0X1C2;
assign {OL1X1C4,OL1X2C3}=OL0X4C3+OL0X3C3+OL0X2C3;
assign {OL1X1C5,OL1X2C4}=OL0X5C4+OL0X4C4+OL0X3C4;
assign {OL1X2C5,OL1X3C4}=OL0X2C4+OL0X1C4;
assign {OL1X1C6,OL1X3C5}=OL0X6C5+OL0X5C5+OL0X4C5;
assign {OL1X2C6,OL1X4C5}=OL0X3C5+OL0X2C5+OL0X1C5;
assign {OL1X1C7,OL1X3C6}=OL0X7C6+OL0X6C6+OL0X5C6;
assign {OL1X2C7,OL1X4C6}=OL0X4C6+OL0X3C6+OL0X2C6;
assign {OL1X1C8,OL1X3C7}=OL0X8C7+OL0X7C7+OL0X6C7;
assign {OL1X2C8,OL1X4C7}=OL0X5C7+OL0X4C7+OL0X3C7;
assign {OL1X3C8,OL1X5C7}=OL0X2C7+OL0X1C7;
assign {OL1X1C9,OL1X4C8}=OL0X9C8+OL0X8C8+OL0X7C8;
assign {OL1X2C9,OL1X5C8}=OL0X6C8+OL0X5C8+OL0X4C8;
assign {OL1X3C9,OL1X6C8}=OL0X3C8+OL0X2C8+OL0X1C8;
assign {OL1X1C10,OL1X4C9}=OL0X10C9+OL0X9C9+OL0X8C9;
assign {OL1X2C10,OL1X5C9}=OL0X7C9+OL0X6C9+OL0X5C9;
assign {OL1X3C10,OL1X6C9}=OL0X4C9+OL0X3C9+OL0X2C9;
assign {OL1X1C11,OL1X4C10}=OL0X11C10+OL0X10C10+OL0X9C10;
assign {OL1X2C11,OL1X5C10}=OL0X8C10+OL0X7C10+OL0X6C10;
assign {OL1X3C11,OL1X6C10}=OL0X5C10+OL0X4C10+OL0X3C10;
assign {OL1X4C11,OL1X7C10}=OL0X2C10+OL0X1C10;
assign {OL1X1C12,OL1X5C11}=OL0X12C11+OL0X11C11+OL0X10C11;
assign {OL1X2C12,OL1X6C11}=OL0X9C11+OL0X8C11+OL0X7C11;
assign {OL1X3C12,OL1X7C11}=OL0X6C11+OL0X5C11+OL0X4C11;
assign {OL1X4C12,OL1X8C11}=OL0X3C11+OL0X2C11+OL0X1C11;
assign {OL1X1C13,OL1X5C12}=OL0X13C12+OL0X12C12+OL0X11C12;
assign {OL1X2C13,OL1X6C12}=OL0X10C12+OL0X9C12+OL0X8C12;
assign {OL1X3C13,OL1X7C12}=OL0X7C12+OL0X6C12+OL0X5C12;
assign {OL1X4C13,OL1X8C12}=OL0X4C12+OL0X3C12+OL0X2C12;
assign {OL1X1C14,OL1X5C13}=OL0X14C13+OL0X13C13+OL0X12C13;
assign {OL1X2C14,OL1X6C13}=OL0X11C13+OL0X10C13+OL0X9C13;
assign {OL1X3C14,OL1X7C13}=OL0X8C13+OL0X7C13+OL0X6C13;
assign {OL1X4C14,OL1X8C13}=OL0X5C13+OL0X4C13+OL0X3C13;
assign {OL1X5C14,OL1X9C13}=OL0X2C13+OL0X1C13;
assign {OL1X1C15,OL1X6C14}=OL0X15C14+OL0X14C14+OL0X13C14;
assign {OL1X2C15,OL1X7C14}=OL0X12C14+OL0X11C14+OL0X10C14;
assign {OL1X3C15,OL1X8C14}=OL0X9C14+OL0X8C14+OL0X7C14;
assign {OL1X4C15,OL1X9C14}=OL0X6C14+OL0X5C14+OL0X4C14;
assign {OL1X5C15,OL1X10C14}=OL0X3C14+OL0X2C14+OL0X1C14;
assign {OL1X1C16,OL1X6C15}=OL0X16C15+OL0X15C15+OL0X14C15;
assign {OL1X2C16,OL1X7C15}=OL0X13C15+OL0X12C15+OL0X11C15;
assign {OL1X3C16,OL1X8C15}=OL0X10C15+OL0X9C15+OL0X8C15;
assign {OL1X4C16,OL1X9C15}=OL0X7C15+OL0X6C15+OL0X5C15;
assign {OL1X5C16,OL1X10C15}=OL0X4C15+OL0X3C15+OL0X2C15;
assign {OL1X1C17,OL1X6C16}=OL0X15C16+OL0X14C16+OL0X13C16;
assign {OL1X2C17,OL1X7C16}=OL0X12C16+OL0X11C16+OL0X10C16;
assign {OL1X3C17,OL1X8C16}=OL0X9C16+OL0X8C16+OL0X7C16;
assign {OL1X4C17,OL1X9C16}=OL0X6C16+OL0X5C16+OL0X4C16;
assign {OL1X5C17,OL1X10C16}=OL0X3C16+OL0X2C16+OL0X1C16;
assign {OL1X1C18,OL1X6C17}=OL0X14C17+OL0X13C17+OL0X12C17;
assign {OL1X2C18,OL1X7C17}=OL0X11C17+OL0X10C17+OL0X9C17;
assign {OL1X3C18,OL1X8C17}=OL0X8C17+OL0X7C17+OL0X6C17;
assign {OL1X4C18,OL1X9C17}=OL0X5C17+OL0X4C17+OL0X3C17;
assign {OL1X5C18,OL1X10C17}=OL0X2C17+OL0X1C17;
assign {OL1X1C19,OL1X6C18}=OL0X13C18+OL0X12C18+OL0X11C18;
assign {OL1X2C19,OL1X7C18}=OL0X10C18+OL0X9C18+OL0X8C18;
assign {OL1X3C19,OL1X8C18}=OL0X7C18+OL0X6C18+OL0X5C18;
assign {OL1X4C19,OL1X9C18}=OL0X4C18+OL0X3C18+OL0X2C18;
assign {OL1X1C20,OL1X5C19}=OL0X12C19+OL0X11C19+OL0X10C19;
assign {OL1X2C20,OL1X6C19}=OL0X9C19+OL0X8C19+OL0X7C19;
assign {OL1X3C20,OL1X7C19}=OL0X6C19+OL0X5C19+OL0X4C19;
assign {OL1X4C20,OL1X8C19}=OL0X3C19+OL0X2C19+OL0X1C19;
assign {OL1X1C21,OL1X5C20}=OL0X11C20+OL0X10C20+OL0X9C20;
assign {OL1X2C21,OL1X6C20}=OL0X8C20+OL0X7C20+OL0X6C20;
assign {OL1X3C21,OL1X7C20}=OL0X5C20+OL0X4C20+OL0X3C20;
assign {OL1X4C21,OL1X8C20}=OL0X2C20+OL0X1C20;
assign {OL1X1C22,OL1X5C21}=OL0X10C21+OL0X9C21+OL0X8C21;
assign {OL1X2C22,OL1X6C21}=OL0X7C21+OL0X6C21+OL0X5C21;
assign {OL1X3C22,OL1X7C21}=OL0X4C21+OL0X3C21+OL0X2C21;
assign {OL1X1C23,OL1X4C22}=OL0X9C22+OL0X8C22+OL0X7C22;
assign {OL1X2C23,OL1X5C22}=OL0X6C22+OL0X5C22+OL0X4C22;
assign {OL1X3C23,OL1X6C22}=OL0X3C22+OL0X2C22+OL0X1C22;
assign {OL1X1C24,OL1X4C23}=OL0X8C23+OL0X7C23+OL0X6C23;
assign {OL1X2C24,OL1X5C23}=OL0X5C23+OL0X4C23+OL0X3C23;
assign {OL1X3C24,OL1X6C23}=OL0X2C23+OL0X1C23;
assign {OL1X1C25,OL1X4C24}=OL0X7C24+OL0X6C24+OL0X5C24;
assign {OL1X2C25,OL1X5C24}=OL0X4C24+OL0X3C24+OL0X2C24;
assign {OL1X1C26,OL1X3C25}=OL0X6C25+OL0X5C25+OL0X4C25;
assign {OL1X2C26,OL1X4C25}=OL0X3C25+OL0X2C25+OL0X1C25;
assign {OL1X1C27,OL1X3C26}=OL0X5C26+OL0X4C26+OL0X3C26;
assign {OL1X2C27,OL1X4C26}=OL0X2C26+OL0X1C26;
assign {OL1X1C28,OL1X3C27}=OL0X4C27+OL0X3C27+OL0X2C27;
assign {OL1X1C29,OL1X2C28}=OL0X3C28+OL0X2C28+OL0X1C28;
assign {OL1X1C30,OL1X2C29}=OL0X2C29+OL0X1C29;
//***********************************Begin of Level 2 ************************************
assign {OL2X1C3,FinalOut[2]}=OL1X2C2+OL1X1C2;
assign {OL2X1C4,OL2X2C3}=OL0X1C3+OL1X2C3+OL1X1C3;
assign {OL2X1C5,OL2X2C4}=OL1X3C4+OL1X2C4+OL1X1C4;
assign {OL2X1C6,OL2X2C5}=OL1X4C5+OL1X3C5+OL1X2C5;
assign {OL2X1C7,OL2X2C6}=OL0X1C6+OL1X4C6+OL1X3C6;
assign {OL2X2C7,OL2X3C6}=OL1X2C6+OL1X1C6;
assign {OL2X1C8,OL2X3C7}=OL1X5C7+OL1X4C7+OL1X3C7;
assign {OL2X2C8,OL2X4C7}=OL1X2C7+OL1X1C7;
assign {OL2X1C9,OL2X3C8}=OL1X6C8+OL1X5C8+OL1X4C8;
assign {OL2X2C9,OL2X4C8}=OL1X3C8+OL1X2C8+OL1X1C8;
assign {OL2X1C10,OL2X3C9}=OL0X1C9+OL1X6C9+OL1X5C9;
assign {OL2X2C10,OL2X4C9}=OL1X4C9+OL1X3C9+OL1X2C9;
assign {OL2X1C11,OL2X3C10}=OL1X7C10+OL1X6C10+OL1X5C10;
assign {OL2X2C11,OL2X4C10}=OL1X4C10+OL1X3C10+OL1X2C10;
assign {OL2X1C12,OL2X3C11}=OL1X8C11+OL1X7C11+OL1X6C11;
assign {OL2X2C12,OL2X4C11}=OL1X5C11+OL1X4C11+OL1X3C11;
assign {OL2X3C12,OL2X5C11}=OL1X2C11+OL1X1C11;
assign {OL2X1C13,OL2X4C12}=OL0X1C12+OL1X8C12+OL1X7C12;
assign {OL2X2C13,OL2X5C12}=OL1X6C12+OL1X5C12+OL1X4C12;
assign {OL2X3C13,OL2X6C12}=OL1X3C12+OL1X2C12+OL1X1C12;
assign {OL2X1C14,OL2X4C13}=OL1X9C13+OL1X8C13+OL1X7C13;
assign {OL2X2C14,OL2X5C13}=OL1X6C13+OL1X5C13+OL1X4C13;
assign {OL2X3C14,OL2X6C13}=OL1X3C13+OL1X2C13+OL1X1C13;
assign {OL2X1C15,OL2X4C14}=OL1X10C14+OL1X9C14+OL1X8C14;
assign {OL2X2C15,OL2X5C14}=OL1X7C14+OL1X6C14+OL1X5C14;
assign {OL2X3C15,OL2X6C14}=OL1X4C14+OL1X3C14+OL1X2C14;
assign {OL2X1C16,OL2X4C15}=OL0X1C15+OL1X10C15+OL1X9C15;
assign {OL2X2C16,OL2X5C15}=OL1X8C15+OL1X7C15+OL1X6C15;
assign {OL2X3C16,OL2X6C15}=OL1X5C15+OL1X4C15+OL1X3C15;
assign {OL2X4C16,OL2X7C15}=OL1X2C15+OL1X1C15;
assign {OL2X1C17,OL2X5C16}=OL1X10C16+OL1X9C16+OL1X8C16;
assign {OL2X2C17,OL2X6C16}=OL1X7C16+OL1X6C16+OL1X5C16;
assign {OL2X3C17,OL2X7C16}=OL1X4C16+OL1X3C16+OL1X2C16;
assign {OL2X1C18,OL2X4C17}=OL1X10C17+OL1X9C17+OL1X8C17;
assign {OL2X2C18,OL2X5C17}=OL1X7C17+OL1X6C17+OL1X5C17;
assign {OL2X3C18,OL2X6C17}=OL1X4C17+OL1X3C17+OL1X2C17;
assign {OL2X1C19,OL2X4C18}=OL0X1C18+OL1X9C18+OL1X8C18;
assign {OL2X2C19,OL2X5C18}=OL1X7C18+OL1X6C18+OL1X5C18;
assign {OL2X3C19,OL2X6C18}=OL1X4C18+OL1X3C18+OL1X2C18;
assign {OL2X1C20,OL2X4C19}=OL1X8C19+OL1X7C19+OL1X6C19;
assign {OL2X2C20,OL2X5C19}=OL1X5C19+OL1X4C19+OL1X3C19;
assign {OL2X3C20,OL2X6C19}=OL1X2C19+OL1X1C19;
assign {OL2X1C21,OL2X4C20}=OL1X8C20+OL1X7C20+OL1X6C20;
assign {OL2X2C21,OL2X5C20}=OL1X5C20+OL1X4C20+OL1X3C20;
assign {OL2X3C21,OL2X6C20}=OL1X2C20+OL1X1C20;
assign {OL2X1C22,OL2X4C21}=OL0X1C21+OL1X7C21+OL1X6C21;
assign {OL2X2C22,OL2X5C21}=OL1X5C21+OL1X4C21+OL1X3C21;
assign {OL2X3C22,OL2X6C21}=OL1X2C21+OL1X1C21;
assign {OL2X1C23,OL2X4C22}=OL1X6C22+OL1X5C22+OL1X4C22;
assign {OL2X2C23,OL2X5C22}=OL1X3C22+OL1X2C22+OL1X1C22;
assign {OL2X1C24,OL2X3C23}=OL1X6C23+OL1X5C23+OL1X4C23;
assign {OL2X2C24,OL2X4C23}=OL1X3C23+OL1X2C23+OL1X1C23;
assign {OL2X1C25,OL2X3C24}=OL0X1C24+OL1X5C24+OL1X4C24;
assign {OL2X2C25,OL2X4C24}=OL1X3C24+OL1X2C24+OL1X1C24;
assign {OL2X1C26,OL2X3C25}=OL1X4C25+OL1X3C25+OL1X2C25;
assign {OL2X1C27,OL2X2C26}=OL1X4C26+OL1X3C26+OL1X2C26;
assign {OL2X1C28,OL2X2C27}=OL0X1C27+OL1X3C27+OL1X2C27;
assign {OL2X1C29,OL2X2C28}=OL1X2C28+OL1X1C28;
assign {OL2X1C30,OL2X2C29}=OL1X2C29+OL1X1C29;
assign {OL2X1C31,OL2X2C30}=OL0X1C30+OL1X1C30;
//***********************************Begin of Level 3 ************************************
assign {OL3X1C4,FinalOut[3]}=OL2X2C3+OL2X1C3;
assign {OL3X1C5,OL3X2C4}=OL2X2C4+OL2X1C4;
assign {OL3X1C6,OL3X2C5}=OL1X1C5+OL2X2C5+OL2X1C5;
assign {OL3X1C7,OL3X2C6}=OL2X3C6+OL2X2C6+OL2X1C6;
assign {OL3X1C8,OL3X2C7}=OL2X4C7+OL2X3C7+OL2X2C7;
assign {OL3X1C9,OL3X2C8}=OL2X4C8+OL2X3C8+OL2X2C8;
assign {OL3X1C10,OL3X2C9}=OL1X1C9+OL2X4C9+OL2X3C9;
assign {OL3X2C10,OL3X3C9}=OL2X2C9+OL2X1C9;
assign {OL3X1C11,OL3X3C10}=OL1X1C10+OL2X4C10+OL2X3C10;
assign {OL3X2C11,OL3X4C10}=OL2X2C10+OL2X1C10;
assign {OL3X1C12,OL3X3C11}=OL2X5C11+OL2X4C11+OL2X3C11;
assign {OL3X2C12,OL3X4C11}=OL2X2C11+OL2X1C11;
assign {OL3X1C13,OL3X3C12}=OL2X6C12+OL2X5C12+OL2X4C12;
assign {OL3X2C13,OL3X4C12}=OL2X3C12+OL2X2C12+OL2X1C12;
assign {OL3X1C14,OL3X3C13}=OL2X6C13+OL2X5C13+OL2X4C13;
assign {OL3X2C14,OL3X4C13}=OL2X3C13+OL2X2C13+OL2X1C13;
assign {OL3X1C15,OL3X3C14}=OL1X1C14+OL2X6C14+OL2X5C14;
assign {OL3X2C15,OL3X4C14}=OL2X4C14+OL2X3C14+OL2X2C14;
assign {OL3X1C16,OL3X3C15}=OL2X7C15+OL2X6C15+OL2X5C15;
assign {OL3X2C16,OL3X4C15}=OL2X4C15+OL2X3C15+OL2X2C15;
assign {OL3X1C17,OL3X3C16}=OL1X1C16+OL2X7C16+OL2X6C16;
assign {OL3X2C17,OL3X4C16}=OL2X5C16+OL2X4C16+OL2X3C16;
assign {OL3X3C17,OL3X5C16}=OL2X2C16+OL2X1C16;
assign {OL3X1C18,OL3X4C17}=OL1X1C17+OL2X6C17+OL2X5C17;
assign {OL3X2C18,OL3X5C17}=OL2X4C17+OL2X3C17+OL2X2C17;
assign {OL3X1C19,OL3X3C18}=OL1X1C18+OL2X6C18+OL2X5C18;
assign {OL3X2C19,OL3X4C18}=OL2X4C18+OL2X3C18+OL2X2C18;
assign {OL3X1C20,OL3X3C19}=OL2X6C19+OL2X5C19+OL2X4C19;
assign {OL3X2C20,OL3X4C19}=OL2X3C19+OL2X2C19+OL2X1C19;
assign {OL3X1C21,OL3X3C20}=OL2X6C20+OL2X5C20+OL2X4C20;
assign {OL3X2C21,OL3X4C20}=OL2X3C20+OL2X2C20+OL2X1C20;
assign {OL3X1C22,OL3X3C21}=OL2X6C21+OL2X5C21+OL2X4C21;
assign {OL3X2C22,OL3X4C21}=OL2X3C21+OL2X2C21+OL2X1C21;
assign {OL3X1C23,OL3X3C22}=OL2X5C22+OL2X4C22+OL2X3C22;
assign {OL3X2C23,OL3X4C22}=OL2X2C22+OL2X1C22;
assign {OL3X1C24,OL3X3C23}=OL2X4C23+OL2X3C23+OL2X2C23;
assign {OL3X1C25,OL3X2C24}=OL2X4C24+OL2X3C24+OL2X2C24;
assign {OL3X1C26,OL3X2C25}=OL1X1C25+OL2X3C25+OL2X2C25;
assign {OL3X1C27,OL3X2C26}=OL1X1C26+OL2X2C26+OL2X1C26;
assign {OL3X1C28,OL3X2C27}=OL1X1C27+OL2X2C27+OL2X1C27;
assign {OL3X1C29,OL3X2C28}=OL2X2C28+OL2X1C28;
assign {OL3X1C30,OL3X2C29}=OL2X2C29+OL2X1C29;
assign {OL3X1C31,OL3X2C30}=OL2X2C30+OL2X1C30;
//***********************************Begin of Level 4 ************************************
assign {OL4X1C5,FinalOut[4]}=OL3X2C4+OL3X1C4;
assign {OL4X1C6,OL4X2C5}=OL3X2C5+OL3X1C5;
assign {OL4X1C7,OL4X2C6}=OL3X2C6+OL3X1C6;
assign {OL4X1C8,OL4X2C7}=OL2X1C7+OL3X2C7+OL3X1C7;
assign {OL4X1C9,OL4X2C8}=OL2X1C8+OL3X2C8+OL3X1C8;
assign {OL4X1C10,OL4X2C9}=OL3X3C9+OL3X2C9+OL3X1C9;
assign {OL4X1C11,OL4X2C10}=OL3X4C10+OL3X3C10+OL3X2C10;
assign {OL4X1C12,OL4X2C11}=OL3X4C11+OL3X3C11+OL3X2C11;
assign {OL4X1C13,OL4X2C12}=OL3X4C12+OL3X3C12+OL3X2C12;
assign {OL4X1C14,OL4X2C13}=OL3X4C13+OL3X3C13+OL3X2C13;
assign {OL4X1C15,OL4X2C14}=OL2X1C14+OL3X4C14+OL3X3C14;
assign {OL4X2C15,OL4X3C14}=OL3X2C14+OL3X1C14;
assign {OL4X1C16,OL4X3C15}=OL2X1C15+OL3X4C15+OL3X3C15;
assign {OL4X2C16,OL4X4C15}=OL3X2C15+OL3X1C15;
assign {OL4X1C17,OL4X3C16}=OL3X5C16+OL3X4C16+OL3X3C16;
assign {OL4X2C17,OL4X4C16}=OL3X2C16+OL3X1C16;
assign {OL4X1C18,OL4X3C17}=OL2X1C17+OL3X5C17+OL3X4C17;
assign {OL4X2C18,OL4X4C17}=OL3X3C17+OL3X2C17+OL3X1C17;
assign {OL4X1C19,OL4X3C18}=OL2X1C18+OL3X4C18+OL3X3C18;
assign {OL4X2C19,OL4X4C18}=OL3X2C18+OL3X1C18;
assign {OL4X1C20,OL4X3C19}=OL3X4C19+OL3X3C19+OL3X2C19;
assign {OL4X1C21,OL4X2C20}=OL3X4C20+OL3X3C20+OL3X2C20;
assign {OL4X1C22,OL4X2C21}=OL3X4C21+OL3X3C21+OL3X2C21;
assign {OL4X1C23,OL4X2C22}=OL3X4C22+OL3X3C22+OL3X2C22;
assign {OL4X1C24,OL4X2C23}=OL2X1C23+OL3X3C23+OL3X2C23;
assign {OL4X1C25,OL4X2C24}=OL2X1C24+OL3X2C24+OL3X1C24;
assign {OL4X1C26,OL4X2C25}=OL2X1C25+OL3X2C25+OL3X1C25;
assign {OL4X1C27,OL4X2C26}=OL3X2C26+OL3X1C26;
assign {OL4X1C28,OL4X2C27}=OL3X2C27+OL3X1C27;
assign {OL4X1C29,OL4X2C28}=OL3X2C28+OL3X1C28;
assign {OL4X1C30,OL4X2C29}=OL3X2C29+OL3X1C29;
assign {OL4X1C31,OL4X2C30}=OL3X2C30+OL3X1C30;
assign {OL4X1C32,OL4X2C31}=OL2X1C31+OL3X1C31;
//***********************************Begin of Level 5 ************************************
assign {OL5X1C6,FinalOut[5]}=OL4X2C5+OL4X1C5;
assign {OL5X1C7,OL5X2C6}=OL4X2C6+OL4X1C6;
assign {OL5X1C8,OL5X2C7}=OL4X2C7+OL4X1C7;
assign {OL5X1C9,OL5X2C8}=OL4X2C8+OL4X1C8;
assign {OL5X1C10,OL5X2C9}=OL4X2C9+OL4X1C9;
assign {OL5X1C11,OL5X2C10}=OL3X1C10+OL4X2C10+OL4X1C10;
assign {OL5X1C12,OL5X2C11}=OL3X1C11+OL4X2C11+OL4X1C11;
assign {OL5X1C13,OL5X2C12}=OL3X1C12+OL4X2C12+OL4X1C12;
assign {OL5X1C14,OL5X2C13}=OL3X1C13+OL4X2C13+OL4X1C13;
assign {OL5X1C15,OL5X2C14}=OL4X3C14+OL4X2C14+OL4X1C14;
assign {OL5X1C16,OL5X2C15}=OL4X4C15+OL4X3C15+OL4X2C15;
assign {OL5X1C17,OL5X2C16}=OL4X4C16+OL4X3C16+OL4X2C16;
assign {OL5X1C18,OL5X2C17}=OL4X4C17+OL4X3C17+OL4X2C17;
assign {OL5X1C19,OL5X2C18}=OL4X4C18+OL4X3C18+OL4X2C18;
assign {OL5X1C20,OL5X2C19}=OL3X1C19+OL4X3C19+OL4X2C19;
assign {OL5X1C21,OL5X2C20}=OL3X1C20+OL4X2C20+OL4X1C20;
assign {OL5X1C22,OL5X2C21}=OL3X1C21+OL4X2C21+OL4X1C21;
assign {OL5X1C23,OL5X2C22}=OL3X1C22+OL4X2C22+OL4X1C22;
assign {OL5X1C24,OL5X2C23}=OL3X1C23+OL4X2C23+OL4X1C23;
assign {OL5X1C25,OL5X2C24}=OL4X2C24+OL4X1C24;
assign {OL5X1C26,OL5X2C25}=OL4X2C25+OL4X1C25;
assign {OL5X1C27,OL5X2C26}=OL4X2C26+OL4X1C26;
assign {OL5X1C28,OL5X2C27}=OL4X2C27+OL4X1C27;
assign {OL5X1C29,OL5X2C28}=OL4X2C28+OL4X1C28;
assign {OL5X1C30,OL5X2C29}=OL4X2C29+OL4X1C29;
assign {OL5X1C31,OL5X2C30}=OL4X2C30+OL4X1C30;
assign {OL5X1C32,OL5X2C31}=OL4X2C31+OL4X1C31;
//***********************************Begin of Level 6 ************************************
assign {OL6X1C7,FinalOut[6]}=OL5X2C6+OL5X1C6;
assign {OL6X1C8,OL6X2C7}=OL5X2C7+OL5X1C7;
assign {OL6X1C9,OL6X2C8}=OL5X2C8+OL5X1C8;
assign {OL6X1C10,OL6X2C9}=OL5X2C9+OL5X1C9;
assign {OL6X1C11,OL6X2C10}=OL5X2C10+OL5X1C10;
assign {OL6X1C12,OL6X2C11}=OL5X2C11+OL5X1C11;
assign {OL6X1C13,OL6X2C12}=OL5X2C12+OL5X1C12;
assign {OL6X1C14,OL6X2C13}=OL5X2C13+OL5X1C13;
assign {OL6X1C15,OL6X2C14}=OL5X2C14+OL5X1C14+carry;
assign {OL6X1C16,OL6X2C15}=OL4X1C15+OL5X2C15+OL5X1C15;
assign {OL6X1C17,OL6X2C16}=OL4X1C16+OL5X2C16+OL5X1C16;
assign {OL6X1C18,OL6X2C17}=OL4X1C17+OL5X2C17+OL5X1C17;
assign {OL6X1C19,OL6X2C18}=OL4X1C18+OL5X2C18+OL5X1C18;
assign {OL6X1C20,OL6X2C19}=OL4X1C19+OL5X2C19+OL5X1C19;
assign {OL6X1C21,OL6X2C20}=OL5X2C20+OL5X1C20;
assign {OL6X1C22,OL6X2C21}=OL5X2C21+OL5X1C21;
assign {OL6X1C23,OL6X2C22}=OL5X2C22+OL5X1C22;
assign {OL6X1C24,OL6X2C23}=OL5X2C23+OL5X1C23;
assign {OL6X1C25,OL6X2C24}=OL5X2C24+OL5X1C24;
assign {OL6X1C26,OL6X2C25}=OL5X2C25+OL5X1C25;
assign {OL6X1C27,OL6X2C26}=OL5X2C26+OL5X1C26;
assign {OL6X1C28,OL6X2C27}=OL5X2C27+OL5X1C27;
assign {OL6X1C29,OL6X2C28}=OL5X2C28+OL5X1C28;
assign {OL6X1C30,OL6X2C29}=OL5X2C29+OL5X1C29;
assign {OL6X1C31,OL6X2C30}=OL5X2C30+OL5X1C30;
assign {OL6X1C32,OL6X2C31}=OL5X2C31+OL5X1C31;
wire [24:0] O1,O2;
assign O1[0]=OL6X1C7;
assign O2[0]=OL6X2C7;
assign O1[1]=OL6X1C8;
assign O2[1]=OL6X2C8;
assign O1[2]=OL6X1C9;
assign O2[2]=OL6X2C9;
assign O1[3]=OL6X1C10;
assign O2[3]=OL6X2C10;
assign O1[4]=OL6X1C11;
assign O2[4]=OL6X2C11;
assign O1[5]=OL6X1C12;
assign O2[5]=OL6X2C12;
assign O1[6]=OL6X1C13;
assign O2[6]=OL6X2C13;
assign O1[7]=OL6X1C14;
assign O2[7]=OL6X2C14;
assign O1[8]=OL6X1C15;
assign O2[8]=OL6X2C15;
assign O1[9]=OL6X1C16;
assign O2[9]=OL6X2C16;
assign O1[10]=OL6X1C17;
assign O2[10]=OL6X2C17;
assign O1[11]=OL6X1C18;
assign O2[11]=OL6X2C18;
assign O1[12]=OL6X1C19;
assign O2[12]=OL6X2C19;
assign O1[13]=OL6X1C20;
assign O2[13]=OL6X2C20;
assign O1[14]=OL6X1C21;
assign O2[14]=OL6X2C21;
assign O1[15]=OL6X1C22;
assign O2[15]=OL6X2C22;
assign O1[16]=OL6X1C23;
assign O2[16]=OL6X2C23;
assign O1[17]=OL6X1C24;
assign O2[17]=OL6X2C24;
assign O1[18]=OL6X1C25;
assign O2[18]=OL6X2C25;
assign O1[19]=OL6X1C26;
assign O2[19]=OL6X2C26;
assign O1[20]=OL6X1C27;
assign O2[20]=OL6X2C27;
assign O1[21]=OL6X1C28;
assign O2[21]=OL6X2C28;
assign O1[22]=OL6X1C29;
assign O2[22]=OL6X2C29;
assign O1[23]=OL6X1C30;
assign O2[23]=OL6X2C30;
assign O1[24]=OL6X1C31;
assign O2[24]=OL6X2C31;
assign FinalOut[31:7]=O1+O2;
assign FinalOut_MSB=FinalOut[31:15];
assign FinalOut_LSB=FinalOut[14:0];
endmodule



module ARTS_n32_ss16(A,B,OUT);
input [31:0]A,B;
output reg[63:0]OUT;
//******************* wires ****************************

	wire Ka,Kb;
	wire [15:0]AH,BH,AL,BL;
	wire [14:0]PP1;
	wire carry;
	wire [16:0]Mult_MSB;
	wire [14:0]Mult_LSB;
	wire [14:0]middle_part;
	wire orout1,orout2,z;

	LSD_n32_ss16  S1 (A,Ka,AH,AL);
	LSD_n32_ss16  S2 (B,Kb,BH,BL);
	APPR  S3 (AH,AL,BH,BL,PP1,carry);
	wallace_with_carry mult1 (AH,BH,carry,Mult_MSB,Mult_LSB);
	assign middle_part= Mult_LSB | PP1;
   	assign orout1=AH[0]|AH[1]|AH[2]|AH[3]|AH[4]|AH[5]|AH[6]|AH[7]|AH[8]|AH[9]|AH[10]|AH[11]|AH[12]|AH[13]|AH[14]|AH[15];
	assign orout2=BH[0]|BH[1]|BH[2]|BH[3]|BH[4]|BH[5]|BH[6]|BH[7]|BH[8]|BH[9]|BH[10]|BH[11]|BH[12]|BH[13]|BH[14]|BH[15];
	assign z= orout1 & orout2;
	wire [1:0] my_case;
	assign my_case = (z == 1'b0) ? 2'd0 :
		((Ka==1'd1 && Kb==1'd1)) ? 2'd1:
		((Ka==1'd1 && Kb==1'd0)||(Ka== 1'd0 && Kb==1'd1)) ? 2'd2:2'd3;
	always@(my_case, Mult_MSB, middle_part)begin
		case (my_case)
		2'd0:OUT = 64'b0 ;
		2'd1:OUT = {Mult_MSB, middle_part,32'd4294967295};
		2'd2:OUT = {16'b0, Mult_MSB, middle_part,16'd65535};
		2'd3:OUT = {32'b0, Mult_MSB, middle_part};
		endcase
	end
endmodule

