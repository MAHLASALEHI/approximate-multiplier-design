// n=16 w=2              


module APPR (AH,AL,BH,BL,PP1,carry);
	input [1:0]AH,BH,AL,BL;
	output PP1;
	output carry;
	wire P6,O6,P7,O7;

	assign P6=(BL[1]&AH[1]);
	assign P7=P6;

	assign O6=(AL[1]&BH[1]);
	assign O7=O6;

	assign PP1=P6|O6;
	assign carry= P7|O7;
endmodule

//******************* LSD ***************************
module LSD_n16_ss2(X,Kx,XH,XL);
	input [15:0]X;
	output [2:0]Kx;
	output [1:0]XH;
	output [1:0]XL;
	assign Kx=(X[15] | X[14]) ? 3'b111:
	(X[13] | X[12]) ? 3'b110:
	(X[11] | X[10]) ? 3'b101:
	(X[9] | X[8]) ? 3'b100:
	(X[7] | X[6]) ? 3'b011:
	(X[5] | X[4]) ? 3'b010:
	(X[3] | X[2]) ? 3'b001: 3'b000;

	assign XH=(Kx==3'b111) ? X[15:14]:
	(Kx==3'b110) ? X[13:12]:
	(Kx==3'b101) ? X[11:10]: 
	(Kx==3'b100) ? X[9:8]:
	(Kx==3'b011) ? X[7:6]:
	(Kx==3'b010) ? X[5:4]:
	(Kx==3'b001) ? X[3:2]:X[1:0];

	assign XL=(Kx==3'b111) ? X[13:12]:
	(Kx==3'b110) ? X[11:10]:
	(Kx==3'b101) ? X[9:8]: 
	(Kx==3'b100) ? X[7:6]:
	(Kx==3'b011) ? X[5:4]:
	(Kx==3'b010) ? X[3:2]:
	(Kx==3'b001) ? X[1:0]:2'b00;
endmodule
//**********************HA and FA***********************
module HA(A,B,sum,carry);
    input A, B;
    output sum, carry;
	assign sum = A ^ B;   // XOR operation for sum
	assign carry = A & B; // AND operation for carry
endmodule


module FA (A,B,cin,sum,cout);
    input A, B, cin;
    output sum, cout;
	assign sum = A ^ B ^ cin;
	assign cout = (A & B) | (cin & (A ^ B));
endmodule

//******************* wallace 4 ***************************
module wallace_with_carry(A,B,carry,FinalOut_MSB,FinalOut_LSB);
input [1:0]A,B;
input carry;
output [2:0]FinalOut_MSB;
output FinalOut_LSB;
wire [3:0] FinalOut;
wire A1B0,A0B1,A2B0,A1B1,A0B2,A3B0,A2B1,A1B2,A0B3,A3B1,A2B2,A1B3,A3B2,A2B3,A3B3;
wire c0;
//**************************************Generating PPs**************
assign FinalOut[0]=A[0] & B[0];
assign A1B0= A[1] & B[0];
assign A0B1= A[0] & B[1];
assign A1B1= A[1] & B[1];

	FA aa0 (A0B1,A1B0,carry,FinalOut[1],c0);
	HA aa1 (A1B1,c0,FinalOut[2],FinalOut[3]);

assign FinalOut_MSB=FinalOut[3:1];
assign FinalOut_LSB=FinalOut[0];
endmodule



module ARTS_n16_ss2(A,B,OUT);
input [15:0]A,B;
output reg[31:0]OUT;
//******************* wires ****************************

	wire [2:0]Ka,Kb;
	wire [1:0]AH,BH,AL,BL;
	wire PP1;
	wire carry;
	wire [2:0]Mult_MSB;
	wire Mult_LSB;
	wire middle_part;
	wire orout1,orout2,z;

	LSD_n16_ss2  S1 (A,Ka,AH,AL);
	LSD_n16_ss2  S2 (B,Kb,BH,BL);
	APPR  S3 (AH,AL,BH,BL,PP1,carry);
	wallace_with_carry mult1 (AH,BH,carry,Mult_MSB,Mult_LSB);
	assign middle_part= Mult_LSB | PP1;
   	assign orout1=AH[0]|AH[1];
	assign orout2=BH[0]|BH[1];
	assign z= orout1 & orout2;
	wire [3:0]my_case;
	assign my_case= (z==1'b0) ? 4'd0:
	     (Ka==3'd7 & Kb==3'd7) ? 4'd1:
		 ((Ka==3'd7 & Kb==3'd6) | (Ka==3'd6 & Kb==3'd7)) ? 4'd2:	 
		 ((Ka==3'd7 & Kb==3'd5) | (Ka==3'd5 & Kb==3'd7) | (Ka==3'd6 & Kb==3'd6)) ? 4'd3:
		 ((Ka==3'd7 & Kb==3'd4) | (Ka==3'd4 & Kb==3'd7) | (Ka==3'd6 & Kb==3'd5) | (Ka==3'd5 & Kb==3'd6)) ? 4'd4:
		 ((Ka==3'd7 & Kb==3'd3) | (Ka==3'd3 & Kb==3'd7) | (Ka==3'd6 & Kb==3'd4) | (Ka==3'd4 & Kb==3'd6) | (Ka==3'd5 & Kb==3'd5)) ? 4'd5:
		 ((Ka==3'd7 & Kb==3'd2) | (Ka==3'd2 & Kb==3'd7) | (Ka==3'd6 & Kb==3'd3) | (Ka==3'd3 & Kb==3'd6) | (Ka==3'd5 & Kb==3'd4) | (Ka==3'd4 & Kb==3'd5)) ? 4'd6:
		 ((Ka==3'd7 & Kb==3'd1) | (Ka==3'd1 & Kb==3'd7) | (Ka==3'd6 & Kb==3'd2) | (Ka==3'd2 & Kb==3'd6) | (Ka==3'd5 & Kb==3'd3) | (Ka==3'd3 & Kb==3'd5) | (Ka==3'd4 & Kb==3'd4)) ? 4'd7:
		 ((Ka==3'd7 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd7) | (Ka==3'd6 & Kb==3'd1) | (Ka==3'd1 & Kb==3'd6) | (Ka==3'd5 & Kb==3'd2) | (Ka==3'd2 & Kb==3'd5) | (Ka==3'd4 & Kb==3'd3) | (Ka==3'd3 & Kb==3'd4)) ? 4'd8:
		 ((Ka==3'd6 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd6) | (Ka==3'd5 & Kb==3'd1) | (Ka==3'd1 & Kb==3'd5) | (Ka==3'd4 & Kb==3'd2) | (Ka==3'd2 & Kb==3'd4) | (Ka==3'd3 & Kb==3'd3)) ? 4'd9:
		 ((Ka==3'd5 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd5) | (Ka==3'd4 & Kb==3'd1) | (Ka==3'd1 & Kb==3'd4) | (Ka==3'd3 & Kb==3'd2) | (Ka==3'd2 & Kb==3'd3)) ? 4'd10:
		 ((Ka==3'd4 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd4) | (Ka==3'd3 & Kb==3'd1) | (Ka==3'd1 & Kb==3'd3) | (Ka==3'd2 & Kb==3'd2)) ? 4'd11:
		 ((Ka==3'd3 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd3) | (Ka==3'd2 & Kb==3'd1) | (Ka==3'd1 & Kb==3'd2)) ? 4'd12:
		 ((Ka==3'd2 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd2) | (Ka==3'd1 & Kb==3'd1)) ? 4'd13:
		 ((Ka==3'd1 & Kb==3'd0) | (Ka==3'd0 & Kb==3'd1)) ? 4'd14: 4'd15;
	always@(my_case, Mult_MSB, middle_part)begin
		case (my_case)
		4'd0: OUT=32'b0;
	    4'd1: OUT={Mult_MSB,middle_part,28'b1111111111111111111111111111} ;
		4'd2: OUT={2'b0,Mult_MSB,middle_part,26'b11111111111111111111111111} ;
		4'd3: OUT={4'b0,Mult_MSB,middle_part,24'b111111111111111111111111} ;
		4'd4: OUT={6'b0,Mult_MSB,middle_part,22'b1111111111111111111111}; 
		4'd5: OUT={8'b0,Mult_MSB,middle_part,20'b11111111111111111111} ;
		4'd6: OUT={10'b0,Mult_MSB,middle_part,18'b111111111111111111} ;
		4'd7: OUT={12'b0,Mult_MSB,middle_part,16'b1111111111111111} ;
		4'd8: OUT={14'b0,Mult_MSB,middle_part,14'b11111111111111} ;
		4'd9: OUT={16'b0,Mult_MSB,middle_part,12'b111111111111};
		4'd10: OUT={18'b0,Mult_MSB,middle_part,10'b1111111111} ;
		4'd11: OUT={20'b0,Mult_MSB,middle_part,8'b11111111} ;
		4'd12: OUT={22'b0,Mult_MSB,middle_part,6'b111111} ;
		4'd13: OUT={24'b0,Mult_MSB,middle_part,4'b1111} ;
		4'd14: OUT={26'b0,Mult_MSB,middle_part,2'b11} ;
		4'd15: OUT={28'd0,Mult_MSB,middle_part};
		endcase
	end
endmodule

